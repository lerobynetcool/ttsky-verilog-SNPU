`default_nettype none

// https://github.com/IHP-GmbH/IHP-Open-PDK/blob/main/ihp-sg13g2/libs.ref/sg13g2_stdcell/verilog/sg13g2_stdcell.v
// type: nand2
`timescale 1ns/10ps
`celldefine
module sg13g2_nand2_1 (Y, A, B);
	output Y;
	input A, B;

	// Function
	wire int_fwire_0;

	and (int_fwire_0, A, B);
	not (Y, int_fwire_0);

	// Timing
	specify
		(A => Y) = 0;
		(B => Y) = 0;
	endspecify
endmodule
`endcelldefine

module nand_latch (
	input wire S,
	input wire R,
	output wire Q,
	output wire Qn
);
	sg13g2_nand2_1 Q_inst (.A(S), .B(Qn), .Y(Q));
	sg13g2_nand2_1 Qn_inst (.A(R), .B(Q), .Y(Qn));
endmodule

module funky_rnd(
	input wire G, // generator state : 0 = random mode, 1 = freeze
	output wire R // output random value between 0 or 1
);
	wire Qn_ignore;
	nand_latch my_latch (
		.S(G), // !!! normally, S=R=0 is banned, but here I want Q to be random
		.R(G), // !!! so it's all good... maybe ? I don't know electronics enough.
		.Q(R),
		.Qn(Qn_ignore)
	);
endmodule
